module MultibitAdder(G11,G12,G14);
input [3:0] G11,G12;
output [3:0]G14;
assign G14=G11+G12;
endmodule
